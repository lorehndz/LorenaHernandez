module Contador 